module memory#(parameter m =32)
				(      input [4:0]PC,
				       output [m-1:0]out
				);	
			reg [m-1:0] Mem [31:0];
			assign out = Mem[PC];
			always@(PC) begin
				Mem[0]= {2'b00,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[1]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[2]= {2'b01,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[3]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[4]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[5]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[6]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[7]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[8]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[9]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[10]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[11]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[12]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[13]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[14]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[15]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[16]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[17]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[18]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[19]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[20]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[21]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[22]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[23]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[24]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[25]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[26]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[27]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[28]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[29]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[30]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				Mem[31]= {2'b10,5'b00100,5'b00101,5'b00000,5'b00001,5'b00010,5'b00011};
				
				
			end		
endmodule
